module microui

import gg

pub fn gg_r_draw_text(ctx &gg.Context, text &char, pos C.mu_Vec2, color C.mu_Color) {
    str := unsafe { cstring_to_vstring(text) }
	// println("draw_text text: ${str}")
	// println("draw_text text: ${text}, pos: ${pos}, color: ${color}")
    ctx.draw_text(pos.x, pos.y, str,
        size:  30
        color: gg.Color{r: color.r, g: color.g, b: color.b, a: color.a}
    )
}

pub fn gg_r_draw_rect(ctx &gg.Context, rect C.mu_Rect, color C.mu_Color) {
    ctx.draw_rect_filled(rect.x, rect.y, rect.w, rect.h, gg.Color{r: color.r, g: color.g, b: color.b, a: color.a})
}

pub fn gg_r_draw_icon(ctx &gg.Context, id i32, rect C.mu_Rect, color C.mu_Color) {
    // workaround
    ctx.draw_rect_filled(rect.x, rect.y, rect.w, rect.h, gg.Color{r: color.r, g: color.g, b: color.b, a: color.a})
}

pub fn gg_r_set_clip_rect(ctx &gg.Context, rect C.mu_Rect) {
    // ctx.set_clip_rect(rect.x, rect.y, rect.w, rect.h)
    // currently do nothing
}

pub fn gg_r_text_width(font C.mu_Font, text &char, len i32) i32 {
  len_ := if len == -1 {
        unsafe { C.strlen(text) }
    }else {
        len
    }
  return unsafe { i32(C.strlen(text)) } // WORKAROUND
//   return r_get_text_width(text, len);
}

pub fn gg_r_text_height(font C.mu_Font) int {
//   return r_get_text_height();
    return 30 // WORKAROUND
}